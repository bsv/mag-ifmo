module fifo
#(
    parameter B = 8, // number of bits in a word
              W = 4  // number of address bits
)
(
    input wire clk, reset,
    input wire rd, wr,
    input wire [B-1:0] w_data,
    output wire empty, full,
    output wire [B-1:0] r_data
);

    reg [B-1:0] array_reg [2**W-1:0];
    reg [W-1:0] w_ptr_reg, w_ptr_next, w_ptr_succ;
    reg [W-1:0] r_ptr_reg, r_ptr_next, r_ptr_succ;
    reg full_reg, empty_reg, full_next, empty_next;
    
    /*initial
    begin
        array_reg[0] = 8'h83;
        array_reg[1] = 8'h55;
        array_reg[2] = 8'h66;
        array_reg[3] = 8'h33;
        array_reg[4] = 8'h22;
        array_reg[5] = 8'h44;
    end*/
    
    wire wr_en;
    
    always @(posedge clk)
        if(wr_en)
            array_reg[w_ptr_reg] <= w_data;
    
    assign r_data = array_reg[r_ptr_reg];
    assign wr_en = wr & ~full_reg;
    assign full = full_reg;
    assign empty = empty_reg;
    
    always@(posedge clk, posedge reset)
        if(reset)
            begin
                w_ptr_reg <= 0;
                r_ptr_reg <= 0;
                full_reg <= 0;
                empty_reg <= 1;
                /*w_ptr_reg <= 6;
                r_ptr_reg <= 0;
                full_reg <= 0;
                empty_reg <= 0;*/
                //==========================
            end
        else
            begin
                w_ptr_reg <= w_ptr_next;
                r_ptr_reg <= r_ptr_next;
                full_reg <= full_next;
                empty_reg <= empty_next;
            end
            
    always@*
    begin
        w_ptr_succ = w_ptr_reg + 1;
        r_ptr_succ = r_ptr_reg + 1;
        w_ptr_next = w_ptr_reg;
        r_ptr_next = r_ptr_reg;
        full_next = full_reg;
        empty_next = empty_reg;
        case({wr, rd})
            // 2'b00 : no op
            2'b01: // read
                if(~empty_reg)
                    begin
                        r_ptr_next = r_ptr_succ;
                        full_next = 0;
                        if(r_ptr_succ == w_ptr_reg)
                            empty_next = 1;
                    end
            2'b10: // write
                if(~full_reg)
                    begin
                        w_ptr_next = w_ptr_succ;
                        empty_next = 0;
                        if(w_ptr_succ == r_ptr_reg)
                            full_next = 1;
                    end
            2'b11: // write and read
                begin
                    w_ptr_next = w_ptr_succ;
                    r_ptr_next = r_ptr_succ;
                end
        endcase
    end

endmodule
